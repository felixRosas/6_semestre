LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY secuencial IS
PORT(
d, clk: 	in std_logic;
Q: 		out std_logic
);
END secuencial;

ARCHITECTURE arqsecuencial OF secuencial IS

BEGIN

PROCESS(clk)
BEGIN
	IF clk = '1' THEN
		Q <= d;
	END IF;
END PROCESS;
			
	
END arqsecuencial;